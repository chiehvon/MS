fdsuhifhalldfaogfuedgou